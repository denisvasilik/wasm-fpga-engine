library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
  use work.WasmFpgaEnginePackage.all;
  use work.WasmFpgaStackWshBn_Package.all;

--
-- end
--
-- A pseudo-instruction that terminates a block.
--
entity InstructionEnd is
    port (
        Clk : in std_logic;
        nRst : in std_logic;
        WasmFpgaInvocation_WasmFpgaInstruction : in T_WasmFpgaInvocation_WasmFpgaInstruction;
        WasmFpgaInstruction_WasmFpgaInvocation : out T_WasmFpgaInstruction_WasmFpgaInvocation;
        WasmFpgaStack_WasmFpgaInstruction : in T_WasmFpgaStack_WasmFpgaInstruction;
        WasmFpgaInstruction_WasmFpgaStack : out T_WasmFpgaInstruction_WasmFpgaStack;
        WasmFpgaModuleRam_WasmFpgaInstruction : in T_WasmFpgaModuleRam_WasmFpgaInstruction;
        WasmFpgaInstruction_WasmFpgaModuleRam : out T_WasmFpgaInstruction_WasmFpgaModuleRam
    );
end entity;

architecture InstructionEndArchitecture of InstructionEnd is

    signal Rst : std_logic;
    signal State : std_logic_vector(15 downto 0);

begin

    Rst <= not nRst;

    -- Stack not used
    WasmFpgaInstruction_WasmFpgaStack.Run <= '0';
    WasmFpgaInstruction_WasmFpgaStack.Action <= '0';
    WasmFpgaInstruction_WasmFpgaStack.TypeValue <= WASMFPGASTACK_VAL_i32;
    WasmFpgaInstruction_WasmFpgaStack.HighValue <= (others => '0');
    WasmFpgaInstruction_WasmFpgaStack.LowValue <= (others => '0');

    -- Module not used
    WasmFpgaInstruction_WasmFpgaModuleRam.Run <= '0';
    WasmFpgaInstruction_WasmFpgaModuleRam.Address <= (others => '0');

    process (Clk, Rst) is
    begin
        if (Rst = '1') then
          WasmFpgaInstruction_WasmFpgaInvocation.Address <= (others => '0');
          WasmFpgaInstruction_WasmFpgaInvocation.Trap <= '0';
          WasmFpgaInstruction_WasmFpgaInvocation.Busy <= '1';
          State <= StateIdle;
        elsif rising_edge(Clk) then
            if (State = StateIdle) then
                WasmFpgaInstruction_WasmFpgaInvocation.Busy <= '0';
                if (WasmFpgaInvocation_WasmFpgaInstruction.Run = '1') then
                    WasmFpgaInstruction_WasmFpgaInvocation.Busy <= '1';
                    WasmFpgaInstruction_WasmFpgaInvocation.Address <= WasmFpgaInvocation_WasmFpgaInstruction.Address;
                    State <= StateIdle;
                end if;
            end if;
        end if;
    end process;

end architecture;